----------------------------------------------------------------------------------
-- Company: Fakulteta za ra�unalni�tvo in informatiko
-- Engineer: Luka Prijatelj
-- Create Date:    19:31:24 01/20/2016 
-- Module Name:    BALL_RAM32x128 - Behavioral  
-- Project Name:		SeminarskaNaloga
-- Target Devices: 	Digilent Nexys 4
-- Tool versions:		ISE Project Suite
-- Description: 
--		Modul, ki se uporablja za branje slik/ikon letal in podobnega.
----------------------------------------------------------------------------------

library IEEE;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;





entity BALL_RAM32x128 is
    Port ( clk_i 		: in  STD_LOGIC;
           addrOUT_i : in  STD_LOGIC_VECTOR (6 downto 0);
           data_o 	: out  STD_LOGIC_VECTOR (0 to 31));
end BALL_RAM32x128;






architecture Behavioral of BALL_RAM32x128 is

	type ram_type is array (127 downto 0) of std_logic_vector (0 to 31);
   signal RAM : ram_type;
	signal dataOUT : STD_LOGIC_VECTOR (0 to 31);

begin

	-- to je dvokanalni RAM. Pisemo na naslov addrIN_i, istocasno lahko beremo z naslova addrOUT_i
	-- RAM ima asinhronski bralni dostop, tako da ga je easy za uporabit. Ko naslovis, takoj dobis podatke.
	-- pisalni dostop je sinhronski.
	-- Pazi LSB bit je skrajno levi, zato da se lazje 'ujema' z organizacijo zaslona!

	data_o <= dataOUT;

	process (clk_i)
	begin
		if (clk_i'event and clk_i = '1') then
			-- ZOGA (Velika)
			RAM(0) <= "00000000000111111111100000000000";
			RAM(1) <= "00000000011111111111111000000000";
			RAM(2) <= "00000001111111111111111110000000";
			RAM(3) <= "00000011111111111111111111000000";
			RAM(4) <= "00000111111111111111111111100000";
			RAM(5) <= "00001111111111111111111111110000";
			RAM(6) <= "00011111111111111111111111111000";
			RAM(7) <= "00111111111111111111111111111100";
			RAM(8) <= "00111111111111111111111111111100";
			RAM(9) <= "01111111111111111111111111111110";
			RAM(10) <= "01111111111111111111111111111110";
			RAM(11) <= "11111111111111111111111111111110";
			RAM(12) <= "11111111111111111111111111111110";
			RAM(13) <= "11111111111111111111111111111111";
			RAM(14) <= "11111111111111111111111111111111";
			RAM(15) <= "11111111111111111111111111111111";
			RAM(16) <= "11111111111111111111111111111111";
			RAM(17) <= "11111111111111111111111111111111";
			RAM(18) <= "11111111111111111111111111111111";
			RAM(19) <= "11111111111111111111111111111111";
			RAM(20) <= "11111111111111111111111111111110";
			RAM(21) <= "01111111111111111111111111111110";
			RAM(22) <= "01111111111111111111111111111110";
			RAM(23) <= "00111111111111111111111111111100";
			RAM(24) <= "00111111111111111111111111111100";
			RAM(25) <= "00011111111111111111111111111000";
			RAM(26) <= "00001111111111111111111111110000";
			RAM(27) <= "00000111111111111111111111100000";
			RAM(28) <= "00000011111111111111111111000000";
			RAM(29) <= "00000001111111111111111110000000";
			RAM(30) <= "00000000011111111111111000000000";
			RAM(31) <= "00000000000111111111100000000000";			

			-- ZOGA (Srednja)
			RAM(32) <= "00000000000000000000000000000000";
			RAM(33) <= "00000000000000000000000000000000";
			RAM(34) <= "00000000000000000000000000000000";
			RAM(35) <= "00000000000000000000000000000000";
			RAM(36) <= "00000000000011111111000000000000";
			RAM(37) <= "00000000001111111111110000000000";
			RAM(38) <= "00000000111111111111111100000000";
			RAM(39) <= "00000001111111111111111110000000";
			RAM(40) <= "00000011111111111111111111000000";
			RAM(41) <= "00000011111111111111111111000000";
			RAM(42) <= "00000111111111111111111111100000";
			RAM(43) <= "00000111111111111111111111100000";
			RAM(44) <= "00001111111111111111111111110000";
			RAM(45) <= "00001111111111111111111111110000";
			RAM(46) <= "00001111111111111111111111110000";
			RAM(47) <= "00001111111111111111111111110000";
			RAM(48) <= "00001111111111111111111111110000";
			RAM(49) <= "00001111111111111111111111110000";
			RAM(50) <= "00001111111111111111111111110000";
			RAM(51) <= "00001111111111111111111111110000";
			RAM(52) <= "00000111111111111111111111100000";
			RAM(53) <= "00000111111111111111111111100000";
			RAM(54) <= "00000011111111111111111111000000";
			RAM(55) <= "00000011111111111111111111000000";
			RAM(56) <= "00000001111111111111111110000000";
			RAM(57) <= "00000000111111111111111100000000";
			RAM(58) <= "00000000001111111111110000000000";
			RAM(59) <= "00000000000011111111000000000000";
			RAM(60) <= "00000000000000000000000000000000";
			RAM(61) <= "00000000000000000000000000000000";
			RAM(62) <= "00000000000000000000000000000000";
			RAM(63) <= "00000000000000000000000000000000";

			-- ZOGA (Mala)
			RAM(64) <= "00000000000000000000000000000000";
			RAM(65) <= "00000000000000000000000000000000";
			RAM(66) <= "00000000000000000000000000000000";
			RAM(67) <= "00000000000000000000000000000000";
			RAM(68) <= "00000000000000000000000000000000";
			RAM(69) <= "00000000000000000000000000000000";
			RAM(70) <= "00000000000000000000000000000000";
			RAM(71) <= "00000000000000000000000000000000";
			RAM(72) <= "00000000000001111110000000000000";
			RAM(73) <= "00000000000111111111100000000000";
			RAM(74) <= "00000000001111111111110000000000";
			RAM(75) <= "00000000011111111111111000000000";
			RAM(76) <= "00000000011111111111111000000000";
			RAM(77) <= "00000000111111111111111100000000";
			RAM(78) <= "00000000111111111111111100000000";
			RAM(79) <= "00000000111111111111111100000000";
			RAM(80) <= "00000000111111111111111100000000";
			RAM(81) <= "00000000111111111111111100000000";
			RAM(82) <= "00000000111111111111111100000000";
			RAM(83) <= "00000000011111111111111000000000";
			RAM(84) <= "00000000011111111111111000000000";
			RAM(85) <= "00000000001111111111110000000000";
			RAM(86) <= "00000000000111111111100000000000";
			RAM(87) <= "00000000000001111110000000000000";
			RAM(88) <= "00000000000000000000000000000000";
			RAM(89) <= "00000000000000000000000000000000";
			RAM(90) <= "00000000000000000000000000000000";
			RAM(91) <= "00000000000000000000000000000000";
			RAM(92) <= "00000000000000000000000000000000";
			RAM(93) <= "00000000000000000000000000000000";
			RAM(94) <= "00000000000000000000000000000000";
			RAM(95) <= "00000000000000000000000000000000";

			-- ZOGA (Zelo majhna)
			RAM(96) <= "00000000000000000000000000000000";
			RAM(97) <= "00000000000000000000000000000000";
			RAM(98) <= "00000000000000000000000000000000";
			RAM(99) <= "00000000000000000000000000000000";
			RAM(100) <= "00000000000000000000000000000000";
			RAM(101) <= "00000000000000000000000000000000";
			RAM(102) <= "00000000000000000000000000000000";
			RAM(103) <= "00000000000000000000000000000000";
			RAM(104) <= "00000000000000000000000000000000";
			RAM(105) <= "00000000000000000000000000000000";
			RAM(106) <= "00000000000000000000000000000000";
			RAM(107) <= "00000000000000000000000000000000";
			RAM(108) <= "00000000000000111100000000000000";
			RAM(109) <= "00000000000001111110000000000000";
			RAM(110) <= "00000000000011111111000000000000";
			RAM(111) <= "00000000000011111111000000000000";
			RAM(112) <= "00000000000011111111000000000000";
			RAM(113) <= "00000000000011111111000000000000";
			RAM(114) <= "00000000000001111110000000000000";
			RAM(115) <= "00000000000000111100000000000000";
			RAM(116) <= "00000000000000000000000000000000";
			RAM(117) <= "00000000000000000000000000000000";
			RAM(118) <= "00000000000000000000000000000000";
			RAM(119) <= "00000000000000000000000000000000";
			RAM(120) <= "00000000000000000000000000000000";
			RAM(121) <= "00000000000000000000000000000000";
			RAM(122) <= "00000000000000000000000000000000";
			RAM(123) <= "00000000000000000000000000000000";
			RAM(124) <= "00000000000000000000000000000000";
			RAM(125) <= "00000000000000000000000000000000";
			RAM(126) <= "00000000000000000000000000000000";
			RAM(127) <= "00000000000000000000000000000000";

			-- 256 = MAX_NUMBER_OF_RAM_LINES_FOR_8_BIT_ADDRESS
		end if;
	end process;

	dataOUT <= RAM(conv_integer(addrOUT_i));

end Behavioral;


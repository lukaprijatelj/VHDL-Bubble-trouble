----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:05:28 08/03/2016 
-- Design Name: 
-- Module Name:    END_SCREEN_RAM80x256 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;




entity END_SCREEN_RAM80x256 is
    Port ( clk_i 		: in  STD_LOGIC;
           addrOUT_i : in  STD_LOGIC_VECTOR (7 downto 0);
           data_o 	: out  STD_LOGIC_VECTOR (0 to 79));
end END_SCREEN_RAM80x256;

architecture Behavioral of END_SCREEN_RAM80x256 is

	type ram_type is array (255 downto 0) of std_logic_vector (0 to 79);
   signal RAM : ram_type;
	signal dataOUT : STD_LOGIC_VECTOR (0 to 79);

begin

	-- to je dvokanalni RAM. Pisemo na naslov addrIN_i, istocasno lahko beremo z naslova addrOUT_i
	-- RAM ima asinhronski bralni dostop, tako da ga je easy za uporabit. Ko naslovis, takoj dobis podatke.
	-- pisalni dostop je sinhronski.
	-- Pazi LSB bit je skrajno levi, zato da se lazje 'ujema' z organizacijo zaslona!

	data_o <= dataOUT;

	process (clk_i)
	begin
		if (clk_i'event and clk_i = '1') then
			-- YOU WON
			RAM(0) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(1) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(2) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(3) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(4) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(5) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(6) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(7) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(8) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(9) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(10) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(11) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(12) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(13) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(14) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(15) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(16) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(17) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(18) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(19) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(20) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(21) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(22) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(23) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(24) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(25) <= "00000000111000111001111100011000011000011100011100011001111100011100001100000000";
			RAM(26) <= "00000000111100111011111110011000011000011100011100111011111110011110001100000000";
			RAM(27) <= "00000000011101110111001111011000011000001100111100111111100111011111001100000000";
			RAM(28) <= "00000000001111100110000111011000011000001100111100110111000011011111001100000000";
			RAM(29) <= "00000000001111101110000011011000011000001110111110110110000011111111101100000000";
			RAM(30) <= "00000000000111001110000011011000011000001110110111110110000011111101101100000000";
			RAM(31) <= "00000000000111001110000111011000011000000111100111110111000011111100111100000000";
			RAM(32) <= "00000000000111000111000111011100111000000111100111100111000111011100111100000000";
			RAM(33) <= "00000000000111000111111110011111111000000111100111100011111111011100011100000000";
			RAM(34) <= "00000000000111000011111100001111110000000011100011100001111110011100001100000000";
			RAM(35) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(36) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(37) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(38) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(39) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(40) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(41) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(42) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(43) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(44) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(45) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(46) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(47) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(48) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(49) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(50) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(51) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(52) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(53) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(54) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(55) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(56) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(57) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(58) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(59) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";

			-- YOU LOST
			RAM(60) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(61) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(62) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(63) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(64) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(65) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(66) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(67) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(68) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(69) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(70) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(71) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(72) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(73) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(74) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(75) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(76) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(77) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(78) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(79) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(80) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(81) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(82) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(83) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(84) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(85) <= "00000000111000111001111100011000011000001100000011111000011111011111111000000000";
			RAM(86) <= "00000000111100111011111110011000011000001100000111111100111111011111111000000000";
			RAM(87) <= "00000000011101110111001111011000011000001100001110001110111000000111000000000000";
			RAM(88) <= "00000000001111100110000111011000011000001100001100000110111000000111000000000000";
			RAM(89) <= "00000000001111101110000011011000011000001100001100000110111110000111000000000000";
			RAM(90) <= "00000000000111001110000011011000011000001100001100000110011111000111000000000000";
			RAM(91) <= "00000000000111001110000111011000011000001100001100000110000111100111000000000000";
			RAM(92) <= "00000000000111000111000111011100111000001100001110001110000011100111000000000000";
			RAM(93) <= "00000000000111000111111110011111111000001111110111111100111111000111000000000000";
			RAM(94) <= "00000000000111000011111100001111110000001111110011111000111111000111000000000000";
			RAM(95) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(96) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(97) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(98) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(99) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(100) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(101) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(102) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(103) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(104) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(105) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(106) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(107) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(108) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(109) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(110) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(111) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(112) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(113) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(114) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(115) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(116) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(117) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(118) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(119) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";

			-- PAUSE
			RAM(120) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(121) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(122) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(123) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(124) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(125) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(126) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(127) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(128) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(129) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(130) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(131) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(132) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(133) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(134) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(135) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(136) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(137) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(138) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(139) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(140) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(141) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(142) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(143) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(144) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(145) <= "00000000000000000000111111000011100001100001100111110111111000000000000000000000";
			RAM(146) <= "00000000000000000000111111100111100001100001101111110111111000000000000000000000";
			RAM(147) <= "00000000000000000000111001110111110001100001101100000111000000000000000000000000";
			RAM(148) <= "00000000000000000000111001111110110001100001101110000111000000000000000000000000";
			RAM(149) <= "00000000000000000000111001101110110001100001101111100111111000000000000000000000";
			RAM(150) <= "00000000000000000000111111101100111001100001100111110111111000000000000000000000";
			RAM(151) <= "00000000000000000000111111001111111001100001100001110111000000000000000000000000";
			RAM(152) <= "00000000000000000000111000011111111101110011100001110111000000000000000000000000";
			RAM(153) <= "00000000000000000000111000011100011101111111101111110111111100000000000000000000";
			RAM(154) <= "00000000000000000000111000111000001100111111001111110111111100000000000000000000";
			RAM(155) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(156) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(157) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(158) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(159) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(160) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(161) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(162) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(163) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(164) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(165) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(166) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(167) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(168) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(169) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(170) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(171) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(172) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(173) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(174) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(175) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(176) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(177) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(178) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			RAM(179) <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000";
			-- 128 = MAX_NUMBER_OF_RAM_LINES_FOR_8_BIT_ADDRESS
		end if;
	end process;

	dataOUT <= RAM(conv_integer(addrOUT_i));


end Behavioral;

